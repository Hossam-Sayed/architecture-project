module BaudRateGenerator  #(
    parameter CLOCK_RATE = 100000000,
    parameter BAUD_RATE = 115200
)(
    input wire clk,     // CPU clock
    input wire osmSel, // Oversampling mode select x13 or x16
    output reg rxClk, // baud rate for rx
    output reg txClk // baud rate for tx
);

parameter MIN_OVERSAMPLING_MODE = 13;
parameter MAX_RATE_RX = CLOCK_RATE / (2 * BAUD_RATE * MIN_OVERSAMPLING_MODE);
parameter MAX_RATE_TX = CLOCK_RATE / (2 * BAUD_RATE);
parameter RX_CNT_WIDTH = $clog2(MAX_RATE_RX);
parameter TX_CNT_WIDTH = $clog2(MAX_RATE_TX);
parameter MAX_RATE_13x = MAX_RATE_TX / 13;
parameter MAX_RATE_16x = MAX_RATE_TX / 16;

reg [RX_CNT_WIDTH - 1:0] rxCounter = 0;
reg [TX_CNT_WIDTH - 1:0] txCounter = 0;

initial begin
    rxClk = 1'b0;
    txClk = 1'b0;
end

always @(posedge clk) begin
    // rx clock
    if ((rxCounter == MAX_RATE_13x[RX_CNT_WIDTH-1:0]) || (osmSel == 0 && rxCounter == MAX_RATE_16x[RX_CNT_WIDTH-1:0])) begin
        rxCounter <= 0;
        rxClk <= ~rxClk;
    end
    else begin
        rxCounter <= rxCounter + 1;
    end
    // tx clock
    if (txCounter == MAX_RATE_TX[TX_CNT_WIDTH-1:0]) begin
        txCounter <= 0;
        txClk <= ~txClk;
    end
    else begin
        txCounter <= txCounter + 1;
    end
end

endmodule




module BaudGenerator_tb();

  reg clk;    
  reg osmSel; 
  wire rxClk; 
  wire txClk; 

  always
    begin
    #10
    clk = ~clk;
    end

 

  initial 
  begin
    clk = 0;osmSel = 0;
    #30000
    osmSel = 1;
    #30000
   $stop;
  end

BaudRateGenerator gen(
    clk,    
    osmSel, 
    rxClk, 
    txClk 
);

 


endmodule
